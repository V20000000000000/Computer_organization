module Multiplicand (
    output [31:0] multiplicand_out,
    input [31:0] multiplicand_in,
    input w_ctrl_Multiplicand,
    input rst
)

endmodule