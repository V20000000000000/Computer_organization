module Divisor (
    output [31:0] reg1_out,
    input [31:0] reg1_in,
    input w_ctrl_reg1,
    input rst
);
    
    assign reg1_out = reg1_in;

endmodule


