module Control (
    output rdy,
    output w_ctrl_Multiplicand,
    output srl_ctrl,
    output [5:0] addu_ctrl,
    output w_ctrl_Product,
    input run,
    input rst,
    input clk,
    input lsb
)