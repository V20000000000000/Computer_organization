module (
    output [63:0] Prod,
    output Rdy,
    input [31:0] Mult,
    input [31:0] Mul,
    input run,
    input rst,
    input clk
);



endmodule